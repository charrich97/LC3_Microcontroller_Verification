//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit enable_execute_t;
typedef bit [5:0] E_Control_t;
typedef bit [15:0] IR_t;
typedef bit [15:0] npc_in_t;
typedef bit bypass_alu_1_t;
typedef bit bypass_alu_2_t;
typedef bit bypass_mem_1_t;
typedef bit bypass_mem_2_t;
typedef bit [15:0] VSR1_t;
typedef bit [15:0] VSR2_t;
typedef bit [1:0] W_Control_in_t;
typedef bit Mem_Control_in_t;
typedef bit [15:0] Mem_Bypass_Val_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

