//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit [15:0] Data_dout_t;
typedef bit complete_data_t;
typedef bit [15:0] Data_din_t;
typedef bit [15:0] Data_addr_t;
typedef bit Data_rd_t;
typedef bit D_macc_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

