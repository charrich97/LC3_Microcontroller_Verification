//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
//    This interface performs the instruction_memory signal driving.  It is
//     accessed by the uvm instruction_memory driver through a virtual interface
//     handle in the instruction_memory configuration.  It drives the singals passed
//     in through the port connection named bus of type instruction_memory_if.
//
//     Input signals from the instruction_memory_if are assigned to an internal input
//     signal with a _i suffix.  The _i signal should be used for sampling.
//
//     The input signal connections are as follows:
//       bus.signal -> signal_i 
//
//     This bfm drives signals with a _o suffix.  These signals
//     are driven onto signals within instruction_memory_if based on INITIATOR/RESPONDER and/or
//     ARBITRATION/GRANT status.  
//
//     The output signal connections are as follows:
//        signal_o -> bus.signal
//
//                                                                                           
//      Interface functions and tasks used by UVM components:
//
//             configure:
//                   This function gets configuration attributes from the
//                   UVM driver to set any required BFM configuration
//                   variables such as 'initiator_responder'.                                       
//                                                                                           
//             initiate_and_get_response:
//                   This task is used to perform signaling activity for initiating
//                   a protocol transfer.  The task initiates the transfer, using
//                   input data from the initiator struct.  Then the task captures
//                   response data, placing the data into the response struct.
//                   The response struct is returned to the driver class.
//
//             respond_and_wait_for_next_transfer:
//                   This task is used to complete a current transfer as a responder
//                   and then wait for the initiator to start the next transfer.
//                   The task uses data in the responder struct to drive protocol
//                   signals to complete the transfer.  The task then waits for 
//                   the next transfer.  Once the next transfer begins, data from
//                   the initiator is placed into the initiator struct and sent
//                   to the responder sequence for processing to determine 
//                   what data to respond with.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
import uvmf_base_pkg_hdl::*;
import instruction_memory_pkg_hdl::*;
`include "src/instruction_memory_macros.svh"

interface instruction_memory_driver_bfm 
  (instruction_memory_if bus);
  // The following pragma and additional ones in-lined further below are for running this BFM on Veloce
  // pragma attribute instruction_memory_driver_bfm partition_interface_xif

`ifndef XRTL
// This code is to aid in debugging parameter mismatches between the BFM and its corresponding agent.
// Enable this debug by setting UVM_VERBOSITY to UVM_DEBUG
// Setting UVM_VERBOSITY to UVM_DEBUG causes all BFM's and all agents to display their parameter settings.
// All of the messages from this feature have a UVM messaging id value of "CFG"
// The transcript or run.log can be parsed to ensure BFM parameter settings match its corresponding agents parameter settings.
import uvm_pkg::*;
`include "uvm_macros.svh"
initial begin : bfm_vs_agent_parameter_debug
  `uvm_info("CFG", 
      $psprintf("The BFM at '%m' has the following parameters: ", ),
      UVM_DEBUG)
end
`endif

  // Config value to determine if this is an initiator or a responder 
  uvmf_initiator_responder_t initiator_responder;
  // Custom configuration variables.  
  // These are set using the configure function which is called during the UVM connect_phase

  tri clock_i;
  tri reset_i;

  // Signal list (all signals are capable of being inputs and outputs for the sake
  // of supporting both INITIATOR and RESPONDER mode operation. Expectation is that 
  // directionality in the config file was from the point-of-view of the INITIATOR

  // INITIATOR mode input signals
  tri [15:0] Instr_dout_i;
  reg [15:0] Instr_dout_o = 'bz;
  tri  complete_instr_i;
  reg  complete_instr_o = 'bz;

  // INITIATOR mode output signals
  tri  instrmem_rd_i;
  reg  instrmem_rd_o = 'bz;
  tri [15:0] PC_i;
  reg [15:0] PC_o = 'bz;
  tri  I_macc_i;
  reg  I_macc_o = 'bz;

  // Bi-directional signals
  

  assign clock_i = bus.clock;
  assign reset_i = bus.reset;

  // These are signals marked as 'input' by the config file, but the signals will be
  // driven by this BFM if put into RESPONDER mode (flipping all signal directions around)
  assign Instr_dout_i = bus.Instr_dout;
  assign bus.Instr_dout = (initiator_responder == RESPONDER) ? Instr_dout_o : 'bz;
  assign complete_instr_i = bus.complete_instr;
  assign bus.complete_instr = (initiator_responder == RESPONDER) ? complete_instr_o : 'bz;


  // These are signals marked as 'output' by the config file, but the outputs will
  // not be driven by this BFM unless placed in INITIATOR mode.
  assign bus.instrmem_rd = (initiator_responder == INITIATOR) ? instrmem_rd_o : 'bz;
  assign instrmem_rd_i = bus.instrmem_rd;
  assign bus.PC = (initiator_responder == INITIATOR) ? PC_o : 'bz;
  assign PC_i = bus.PC;
  assign bus.I_macc = (initiator_responder == INITIATOR) ? I_macc_o : 'bz;
  assign I_macc_i = bus.I_macc;

  // Proxy handle to UVM driver
  instruction_memory_pkg::instruction_memory_driver   proxy;
  // pragma tbx oneway proxy.my_function_name_in_uvm_driver                 

  // ****************************************************************************
  // **************************************************************************** 
  // Macros that define structs located in instruction_memory_macros.svh
  // ****************************************************************************
  // Struct for passing configuration data from instruction_memory_driver to this BFM
  // ****************************************************************************
  `instruction_memory_CONFIGURATION_STRUCT
  // ****************************************************************************
  // Structs for INITIATOR and RESPONDER data flow
  //*******************************************************************
  // Initiator macro used by instruction_memory_driver and instruction_memory_driver_bfm
  // to communicate initiator driven data to instruction_memory_driver_bfm.           
  `instruction_memory_INITIATOR_STRUCT
    instruction_memory_initiator_s initiator_struct;
  // Responder macro used by instruction_memory_driver and instruction_memory_driver_bfm
  // to communicate Responder driven data to instruction_memory_driver_bfm.
  `instruction_memory_RESPONDER_STRUCT
    instruction_memory_responder_s responder_struct;

  // ****************************************************************************
// pragma uvmf custom reset_condition_and_response begin
  // Always block used to return signals to reset value upon assertion of reset
  always @( posedge reset_i )
     begin
       // RESPONDER mode output signals
       Instr_dout_o <= 'bz;
       complete_instr_o <= 'bz;
       // INITIATOR mode output signals
       instrmem_rd_o <= 'bz;
       PC_o <= 'bz;
       I_macc_o <= 'bz;
       // Bi-directional signals
 
     end    
// pragma uvmf custom reset_condition_and_response end

  // pragma uvmf custom interface_item_additional begin
  // pragma uvmf custom interface_item_additional end

  //******************************************************************
  // The configure() function is used to pass agent configuration
  // variables to the driver BFM.  It is called by the driver within
  // the agent at the beginning of the simulation.  It may be called 
  // during the simulation if agent configuration variables are updated
  // and the driver BFM needs to be aware of the new configuration 
  // variables.
  //

  function void configure(instruction_memory_configuration_s instruction_memory_configuration_arg); // pragma tbx xtf  
    initiator_responder = instruction_memory_configuration_arg.initiator_responder;
  // pragma uvmf custom configure begin
  // pragma uvmf custom configure end
  endfunction                                                                             

// pragma uvmf custom initiate_and_get_response begin
// ****************************************************************************
// UVMF_CHANGE_ME
// This task is used by an initator.  The task first initiates a transfer then
// waits for the responder to complete the transfer.
    task initiate_and_get_response( 
       // This argument passes transaction variables used by an initiator
       // to perform the initial part of a protocol transfer.  The values
       // come from a sequence item created in a sequence.
       input instruction_memory_initiator_s instruction_memory_initiator_struct, 
       // This argument is used to send data received from the responder
       // back to the sequence item.  The sequence item is returned to the sequence.
       output instruction_memory_responder_s instruction_memory_responder_struct 
       );// pragma tbx xtf  
       // 
       // Members within the instruction_memory_initiator_struct:
       //   op_t opcode ;
       //   reg_t sr1 ;
       //   reg_t sr2 ;
       //   reg_t dr ;
       //   im_t im ;
       //   baser_t baser ;
       //   pcoffset9_t pcoffset9 ;
       //   pcoffset6_t pcoffset6 ;
       //   imm5_t imm5 ;
       //   nzp_t nzp ;
       //   bit [15:0] instruction ;
       //   bit complete_instr ;
       //   instrmem_rd_t instrmem_rd ;
       //   bit [16:0] PC ;
       //   bit I_macc ;
       // Members within the instruction_memory_responder_struct:
       //   op_t opcode ;
       //   reg_t sr1 ;
       //   reg_t sr2 ;
       //   reg_t dr ;
       //   im_t im ;
       //   baser_t baser ;
       //   pcoffset9_t pcoffset9 ;
       //   pcoffset6_t pcoffset6 ;
       //   imm5_t imm5 ;
       //   nzp_t nzp ;
       //   bit [15:0] instruction ;
       //   bit complete_instr ;
       //   instrmem_rd_t instrmem_rd ;
       //   bit [16:0] PC ;
       //   bit I_macc ;
       initiator_struct = instruction_memory_initiator_struct;
       //
       // Reference code;
       //    How to wait for signal value
       //      while (control_signal == 1'b1) @(posedge clock_i);
       //    
       //    How to assign a responder struct member, named xyz, from a signal.   
       //    All available initiator input and inout signals listed.
       //    Initiator input signals
       //      instruction_memory_responder_struct.xyz = Instr_dout_i;  //    [15:0] 
       //      instruction_memory_responder_struct.xyz = complete_instr_i;  //     
       //    Initiator inout signals
       //    How to assign a signal from an initiator struct member named xyz.   
       //    All available initiator output and inout signals listed.
       //    Notice the _o.  Those are storage variables that allow for procedural assignment.
       //    Initiator output signals
       //      instrmem_rd_o <= instruction_memory_initiator_struct.xyz;  //     
       //      PC_o <= instruction_memory_initiator_struct.xyz;  //    [15:0] 
       //      I_macc_o <= instruction_memory_initiator_struct.xyz;  //     
       //    Initiator inout signals
    // Initiate a transfer using the data received.
    @(posedge clock_i);
    @(posedge clock_i);
    // Wait for the responder to complete the transfer then place the responder data into 
    // instruction_memory_responder_struct.
    @(posedge clock_i);
    @(posedge clock_i);
    responder_struct = instruction_memory_responder_struct;
  endtask        
// pragma uvmf custom initiate_and_get_response end

// pragma uvmf custom respond_and_wait_for_next_transfer begin
// ****************************************************************************
// The first_transfer variable is used to prevent completing a transfer in the 
// first call to this task.  For the first call to this task, there is not
// current transfer to complete.
bit first_transfer=1;

// UVMF_CHANGE_ME
// This task is used by a responder.  The task first completes the current 
// transfer in progress then waits for the initiator to start the next transfer.
  task respond_and_wait_for_next_transfer( 
       // This argument is used to send data received from the initiator
       // back to the sequence item.  The sequence determines how to respond.
       output instruction_memory_initiator_s instruction_memory_initiator_struct, 
       // This argument passes transaction variables used by a responder
       // to complete a protocol transfer.  The values come from a sequence item.       
       input instruction_memory_responder_s instruction_memory_responder_struct 
       );// pragma tbx xtf   
  // Variables within the instruction_memory_initiator_struct:
  //   op_t opcode ;
  //   reg_t sr1 ;
  //   reg_t sr2 ;
  //   reg_t dr ;
  //   im_t im ;
  //   baser_t baser ;
  //   pcoffset9_t pcoffset9 ;
  //   pcoffset6_t pcoffset6 ;
  //   imm5_t imm5 ;
  //   nzp_t nzp ;
  //   bit [15:0] instruction ;
  //   bit complete_instr ;
  //   instrmem_rd_t instrmem_rd ;
  //   bit [16:0] PC ;
  //   bit I_macc ;
  // Variables within the instruction_memory_responder_struct:
  //   op_t opcode ;
  //   reg_t sr1 ;
  //   reg_t sr2 ;
  //   reg_t dr ;
  //   im_t im ;
  //   baser_t baser ;
  //   pcoffset9_t pcoffset9 ;
  //   pcoffset6_t pcoffset6 ;
  //   imm5_t imm5 ;
  //   nzp_t nzp ;
  //   bit [15:0] instruction ;
  //   bit complete_instr ;
  //   instrmem_rd_t instrmem_rd ;
  //   bit [16:0] PC ;
  //   bit I_macc ;
       // Reference code;
       //    How to wait for signal value
       //      while (control_signal == 1'b1) @(posedge clock_i);
       //    
       //    How to assign a responder struct member, named xyz, from a signal.   
       //    All available responder input and inout signals listed.
       //    Responder input signals
       //      instruction_memory_responder_struct.xyz = instrmem_rd_i;  //     
       //      instruction_memory_responder_struct.xyz = PC_i;  //    [15:0] 
       //      instruction_memory_responder_struct.xyz = I_macc_i;  //     
       //    Responder inout signals
       //    How to assign a signal, named xyz, from an initiator struct member.   
       //    All available responder output and inout signals listed.
       //    Notice the _o.  Those are storage variables that allow for procedural assignment.
       //    Responder output signals
       //      Instr_dout_o <= instruction_memory_initiator_struct.xyz;  //    [15:0] 
       //      complete_instr_o <= instruction_memory_initiator_struct.xyz;  //     
       //    Responder inout signals
  wait(reset_i === 0);
  @(posedge clock_i);
  if(!first_transfer) begin
      Instr_dout_o = instruction_memory_responder_struct.instruction;
      #1 complete_instr_o = instrmem_rd_i;
      @(posedge clock_i);
      #1 complete_instr_o = instrmem_rd_i;
  end
  else begin
    first_transfer= 0;
    Instr_dout_o = instruction_memory_responder_struct.instruction;
    complete_instr_o = instruction_memory_responder_struct.complete_instr;
    @(posedge clock_i);
    complete_instr_o =0;
  end
  endtask
// pragma uvmf custom respond_and_wait_for_next_transfer end

 
endinterface

// pragma uvmf custom external begin
// pragma uvmf custom external end

