//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit [1:0] mem_state_t;
typedef bit M_control_t;
typedef bit [15:0] M_Data_t;
typedef bit [15:0] M_addr_t;
typedef bit [15:0] DMem_dout_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

